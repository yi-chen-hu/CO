module Mux3to1( data0_i, data1_i, data2_i, select_i, data_o );

parameter size = 16;			   
			
//I/O ports               
input wire	[size-1:0] data0_i;          
input wire	[size-1:0] data1_i;
input wire	[size-1:0] data2_i;
input wire	[2-1:0] select_i;
output wire	[size-1:0] data_o; 

//Main function
/*your code here*/

reg [size-1:0] out;
always@(*)
    case(select_i)
        2'b00:  out = data0_i;
        2'b01:  out = data1_i;
        2'b10:  out = data2_i;
        default:out = data0_i;
     endcase

assign data_o = out;

endmodule      
